module example();
myid1
\myid2
myid1
\myid2
endmodule